architecture beh of lab1 is
begin
	Y <= A and (B or C) and (not D);
end beh;